`default_nettype none

module icache_fake (

);

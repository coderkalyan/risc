`default_nettype none

module rob #(
    parameter LEN = 16
) (
    input wire i_clk,
    input wire i_rst_n
);
    
endmodule

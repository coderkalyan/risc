`default_nettype none

module priority_encoder_6bit (
    input wire [63:0] i_vec,
    output reg [5:0] o_code
);
    always @(*) begin
    o_code = 6'h0;

        if (i_vec[0])
            o_code = 6'h0;
        else if (i_vec[1])
            o_code = 6'h1;
        else if (i_vec[2])
            o_code = 6'h2;
        else if (i_vec[3])
            o_code = 6'h3;
        else if (i_vec[4])
            o_code = 6'h4;
        else if (i_vec[5])
            o_code = 6'h5;
        else if (i_vec[6])
            o_code = 6'h6;
        else if (i_vec[7])
            o_code = 6'h7;
        else if (i_vec[8])
            o_code = 6'h8;
        else if (i_vec[9])
            o_code = 6'h9;
        else if (i_vec[10])
            o_code = 6'ha;
        else if (i_vec[11])
            o_code = 6'hb;
        else if (i_vec[12])
            o_code = 6'hc;
        else if (i_vec[13])
            o_code = 6'hd;
        else if (i_vec[14])
            o_code = 6'he;
        else if (i_vec[15])
            o_code = 6'hf;
        else if (i_vec[16])
            o_code = 6'h10;
        else if (i_vec[17])
            o_code = 6'h11;
        else if (i_vec[18])
            o_code = 6'h12;
        else if (i_vec[19])
            o_code = 6'h13;
        else if (i_vec[20])
            o_code = 6'h14;
        else if (i_vec[21])
            o_code = 6'h15;
        else if (i_vec[22])
            o_code = 6'h16;
        else if (i_vec[23])
            o_code = 6'h17;
        else if (i_vec[24])
            o_code = 6'h18;
        else if (i_vec[25])
            o_code = 6'h19;
        else if (i_vec[26])
            o_code = 6'h1a;
        else if (i_vec[27])
            o_code = 6'h1b;
        else if (i_vec[28])
            o_code = 6'h1c;
        else if (i_vec[29])
            o_code = 6'h1d;
        else if (i_vec[30])
            o_code = 6'h1e;
        else if (i_vec[31])
            o_code = 6'h1f;
        else if (i_vec[32])
            o_code = 6'h20;
        else if (i_vec[33])
            o_code = 6'h21;
        else if (i_vec[34])
            o_code = 6'h22;
        else if (i_vec[35])
            o_code = 6'h23;
        else if (i_vec[36])
            o_code = 6'h24;
        else if (i_vec[37])
            o_code = 6'h25;
        else if (i_vec[38])
            o_code = 6'h26;
        else if (i_vec[39])
            o_code = 6'h27;
        else if (i_vec[40])
            o_code = 6'h28;
        else if (i_vec[41])
            o_code = 6'h29;
        else if (i_vec[42])
            o_code = 6'h2a;
        else if (i_vec[43])
            o_code = 6'h2b;
        else if (i_vec[44])
            o_code = 6'h2c;
        else if (i_vec[45])
            o_code = 6'h2d;
        else if (i_vec[46])
            o_code = 6'h2e;
        else if (i_vec[47])
            o_code = 6'h2f;
        else if (i_vec[48])
            o_code = 6'h30;
        else if (i_vec[49])
            o_code = 6'h31;
        else if (i_vec[50])
            o_code = 6'h32;
        else if (i_vec[51])
            o_code = 6'h33;
        else if (i_vec[52])
            o_code = 6'h34;
        else if (i_vec[53])
            o_code = 6'h35;
        else if (i_vec[54])
            o_code = 6'h36;
        else if (i_vec[55])
            o_code = 6'h37;
        else if (i_vec[56])
            o_code = 6'h38;
        else if (i_vec[57])
            o_code = 6'h39;
        else if (i_vec[58])
            o_code = 6'h3a;
        else if (i_vec[59])
            o_code = 6'h3b;
        else if (i_vec[60])
            o_code = 6'h3c;
        else if (i_vec[61])
            o_code = 6'h3d;
        else if (i_vec[62])
            o_code = 6'h3e;
        else if (i_vec[63])
            o_code = 6'h3f;
    end
endmodule
